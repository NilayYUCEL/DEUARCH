ADD_SUB_inst : ADD_SUB PORT MAP (
		add_sub	 => add_sub_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
